LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY halfSplitter IS
  PORT(DIN: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    DOUT: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END halfSplitter;

ARCHITECTURE pchs OF halfSplitter IS
BEGIN
  DOUT <= DIN(31 DOWNTO 16);
END pchs;