LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY memToRegMux IS
  PORT(R0, R1, JAL: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    MEMTOREG, LINK: IN STD_LOGIC;
    ROUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END memToRegMux;

ARCHITECTURE pcMemToRegMux OF memToRegMux IS
BEGIN
  ROUT <= JAL WHEN LINK = '1' ELSE
          R1 WHEN MEMTOREG = '1' ELSE
          R0;
END pcMemToRegMux;