LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY zeroGen IS
  PORT(TOUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END zeroGen;

ARCHITECTURE pczg OF zeroGen IS
BEGIN
  TOUT <= x"00000000";
END pczg;