LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY extender IS
  PORT(PIN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    EXTENDSIGN: IN STD_LOGIC;
    POUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END extender;

ARCHITECTURE pcExtender OF extender IS
BEGIN
  POUT <= x"FFFF" & PIN WHEN PIN(15) = '1' AND EXTENDSIGN = '1' ELSE
         x"0000" & PIN;
END pcExtender;