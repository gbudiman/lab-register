LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY aluctl IS
  PORT(INST: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    ALUOP: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    ACS: OUT STD_LOGIC_VECTOR(2 DOWNTO 0))
END aluctl;

ARCHITECTURE pcaluctl OF aluctl IS
BEGIN
  
END pcaluctl;