LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY splitter IS
  PORT(Q: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    D31_26: OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    D25_21: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    D20_16: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    D15_11: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    D15_0: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    D5_0: OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    D25_0: OUT STD_LOGIC_VECTOR(25 DOWNTO 0));
END splitter;

ARCHITECTURE pcs OF splitter IS
BEGIN
  D31_26 <= Q(31 DOWNTO 26);
  D25_21 <= Q(25 DOWNTO 21);
  D20_16 <= Q(20 DOWNTO 16);
  D15_11 <= Q(15 DOWNTO 11);
  D15_0 <= Q(15 DOWNTO 0);
  D5_0 <= Q(5 DOWNTO 0);
  D25_0 <= Q(25 DOWNTO 0);
END pcs;