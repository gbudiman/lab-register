LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY loadUpperMux IS
  PORT(Q: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    W: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    UPPER: IN STD_LOGIC;
    QOUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END loadUpperMux;

ARCHITECTURE pclum OF loadUpperMux IS
BEGIN
  QOUT <= Q & x"0000" WHEN UPPER = '1' ELSE W;
END pclum;