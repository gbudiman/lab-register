LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY aluSrcMux IS
  PORT(R0: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    R1: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    ALUSRC: IN STD_LOGIC;
    ROUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END aluSrcMux;

ARCHITECTURE pcAluSrcMux OF aluSrcMux IS
BEGIN
  ROUT <= R0 WHEN ALUSRC = '0' ELSE R1;
END pcAluSrcMux;