LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY memToRegMux IS
  PORT(R0: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    R1: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    MEMTOREG: IN STD_LOGIC;
    ROUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END memToRegMux;

ARCHITECTURE pcMemToRegMux OF memToRegMux IS
BEGIN
  ROUT <= R0 WHEN MEMTOREG = '1' ELSE R1;
END pcMemToRegMux;