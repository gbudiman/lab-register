LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY setWriteMux IS
  PORT(ALU, SLT: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    CONTROL: IN STD_LOGIC;
    D: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END setWriteMux;

ARCHITECTURE pcswm OF setWriteMux IS
BEGIN
  D <= SLT WHEN CONTROL = '1' ELSE ALU;
END pcswm;