LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY regMux IS
  PORT(R0: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    R1: IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    REGDST, LINK: IN STD_LOGIC;
    ROUT: OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END regMux;

ARCHITECTURE pcRegMux OF regMux IS
BEGIN
  ROUT <= "11111" WHEN LINK = '1' ELSE
          R1 WHEN REGDST = '1' ELSE
          R0;
END pcRegMux;