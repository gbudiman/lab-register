LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY signExtend IS
  PORT(PIN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    POUT: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END signExtend;

ARCHITECTURE pcSignExtend OF signExtend IS
BEGIN
  POUT <= x"FFFF" & PIN WHEN PIN(15) = '1' ELSE
         x"0000" & PIN;
END pcSignExtend;