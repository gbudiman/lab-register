LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY clu IS
  PORT(QIN: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    LCTL: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    REGDST, EXTSIGN, MEMTOREG, ALUSRC, REGWRITE, MEMWRITE, HALT: OUT STD_LOGIC;
    JREG, JUMP, LINK, BEQ, BNE, SETU, UPPER: OUT STD_LOGIC;
    ALUCTL: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END CLU;

ARCHITECTURE pcclu OF clu IS
  TYPE decodedOperation IS (oADDU, oAND, oJR, oNOR, oOR, oSLT, oSLTU, oSLL, oSRL, oSUBU, oXOR,
    oADDIU, oANDI, oBEQ, oBNE, oLUI, oLW, oORI, oSLTI, oSLTIU, oSW, oXORI, oJ, oJAL, oHALT, oX);
  SIGNAL dcOp: decodedOperation;
BEGIN
  dcOp <= oADDU   WHEN QIN = "000000" AND LCTL = "100001" ELSE -- ADDU
          oAND    WHEN QIN = "000000" AND LCTL = "100100" ELSE -- AND
          oJR     WHEN QIN = "000000" AND LCTL = "001000" ELSE -- JR
          oNOR    WHEN QIN = "000000" AND LCTL = "100111" ELSE -- NOR
          oOR     WHEN QIN = "000000" AND LCTL = "100101" ELSE -- OR
          oSLT    WHEN QIN = "000000" AND LCTL = "101010" ELSE -- SLT
          oSLTU   WHEN QIN = "000000" AND LCTL = "101011" ELSE -- SLTU
          oSLL    WHEN QIN = "000000" AND LCTL = "000000" ELSE -- SLL
          oSRL    WHEN QIN = "000000" AND LCTL = "000010" ELSE -- SRL
          oSUBU   WHEN QIN = "000000" AND LCTL = "100011" ELSE -- SUBU
          oXOR    WHEN QIN = "000000" AND LCTL = "100110" ELSE -- XOR
          
          oADDIU  WHEN QIN = "001001" ELSE -- ADDIU
          oANDI   WHEN QIN = "001100" ELSE -- ANDI
          oBEQ    WHEN QIN = "000100" ELSE -- BEQ
          oBNE    WHEN QIN = "000101" ELSE -- BNE
          oLUI    WHEN QIN = "001111" ELSE -- LUI
          oLW     WHEN QIN = "100011" ELSE -- LW
          oORI    WHEN QIN = "001101" ELSE -- ORI
          oSLTI   WHEN QIN = "001010" ELSE -- SLTI
          oSLTIU  WHEN QIN = "001011" ELSE -- SLTIU
          oSW     WHEN QIN = "101011" ELSE -- SW
          oXORI   WHEN QIN = "001110" ELSE -- XORI
          oJ      WHEN QIN = "000010" ELSE -- J
          oJAL    WHEN QIN = "000011" ELSE -- JAL
          oHALT   WHEN QIN = "111111" ELSE -- HALT
          oX; -- NOP or UNRECOGNIZED OPERATION
END PCCLU;