LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY branchMux IS
  PORT(BEQ, BNE, ZERO: IN STD_LOGIC;
    BRANCHDECS: OUT STD_LOGIC);
END branchMux;

ARCHITECTURE pcbm OF branchMux IS
BEGIN
  BRANCHDECS <= '1' WHEN (BEQ = '1' AND ZERO = '1') OR (BNE = '1' AND ZERO = '0') ELSE '0';
END pcbm;